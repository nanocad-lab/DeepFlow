MACRO system
	package0
	package1
	package2
	package3
	wire(package0, package1)
	wire(package0, package2)
	wire(package0, package3)
	wire(package1, package2)
	wire(package1, package3)
	wire(package2, package3)
END system

MACRO package
	node0
	node1
	node2
	node3
	node4
	node5
	node6
	node7
	write(node0, node1)
	write(node0, node2)
	write(node0, node3)
	write(node1, node2)
	write(node1, node3)
	write(node2, node3)
END package

MACRO node
	accelerator_die
	hbm0
	wire(accelerator_die, hbm0)
	hbm1
	wire(accelerator_die, hbm1)
	hbm2
	wire(accelerator_die, hbm2)
	hbm3
	wire(accelerator_die, hbm3)
END node

MACRO accelerator_die
	network_io0
	network_io1
	network_io2
	network_io3
	noc
	sm0
	sm1
	sm2
	sm3
	mc_phy0
	mc_phy1
	mc_phy2
	mc_phy3
END accelerator_die

MACRO noc
	l2
END noc

MACRO sm
	reg
	core_group
	l1
	wire(reg, core_group)
	wire(core_group, l1)
END sm

MACRO core_group
	core0
	core1
	core2
	core3
END core_group

